// Code your testbench here
// or browse Examples
//`include "RegMem_tb.v"
`include "tb_simple_CPU.v"