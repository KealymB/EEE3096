// Code your design here
`include "alu.v"
`include "CU.v"
`include "RegMem.v"
`include "top.v"